module shifter();